module mod12_counter(
    input clk,
    input reset,
    input enable,
    output reg [3:0] count
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        count <= 4'b0000;
    end
    else if (enable) begin
        if (count == 4'b1011) begin
            count <= 4'b0000;
        end
        else begin
            count <= count + 1'b1;
        end
    end
end

endmodule